HICUM/L2 Output Characteristics Xyce Simulation
.options nonlin reltol=1e-6 abstol=1e-12
.options device temp=26.85

* Netlist
.INCLUDE "bsimsoi_verilog_a.lib"
Ybsimsoi450 M_H n_D n_G 0 0 _0

.PARAM V_G=0
.PARAM V_D=0

VV_G n_G 0 DC {V_G} 
VV_D n_D 0 DC {V_D}

.DC V_D 0 2 0.001 V_G 0.5 0.8 0.01 



.END
