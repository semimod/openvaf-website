Cir

.options reltol=1e-6 vabstol=1e-6 iabstol=1e-12 temp=26.85 save=nooutput

simulator lang = spectre

; Netlist

model bsim bsimbulk type=n version=106.2 \
 LLONG =2E-06 \
 WWIDE =1E-05 \
 TYPE =1 \
 GEOMOD =0 \
 RGEOMOD =0 \
 COVMOD =1 \
 RDSMOD =2 \
 XL =-1.7E-08 \
 XW =1.1E-08 \
 LINT =0 \
 WINT =0 \
 DLC =0 \
 DWC =0 \
 TOXE =1.74E-09 \
 TOXP =1.7E-09 \
 NDEP =4.6E+23 \
 NSD =1E+26 \
 NGATE =8.5E+25 \
 VFB =-1.02 \
 EPSROX =3.9 \
 EPSRSUB =11.9 \
 NI0SUB =1.1E+16 \
 XJ =1.5E-07 \
 DMCG =0 \
 DMDG =0 \
 DMCGT =0 \
 CIT =1E-08 \
 CDSCD =0.001 \
 CDSCB =0 \
 CDSCBL =0.007 \
 CDSCBLEXP =1 \
 NFACTOR =0.002 \
 NFACTORL =2.1E-08 \
 NFACTORLEXP =6.264 \
 NDEPL1 =0.096 \
 NDEPLEXP1 =1 \
 NDEPL2 =-0.0032 \
 NDEPLEXP2 =2.05 \
 DVTP0 =7.5E-07 \
 DVTP1 =-4.4E-07 \
 NDEPW =-0.1548 \
 NDEPWEXP =0.7441 \
 NDEPWL =0 \
 NDEPWLEXP =0.2 \
 K2W =0 \
 GIDLMOD =1 \
 AGIDL =3.728E-08 \
 AGIDLL =-0.04815 \
 AGIDLW =-0.0341 \
 BGIDL =8.123E+09 \
 CGIDL =1.21E-06 \
 EGIDL =-2.952 \
 PHIN =0.05 \
 K2L =0.001636 \
 K2 =-0.014 \
 ETA0 =8.416E-06 \
 ETAB =-5.561E-05 \
 ETABEXP =2.155 \
 DSUB =3 \
 VSAT =6.4E+04 \
 VSATW =0.05 \
 VSATWEXP =1 \
 DELTA =0.15 \
 DELTAL =0.1 \
 DELTALEXP =1E-05 \
 U0 =0.04546 \
 ETAMOB =1.5 \
 U0L =0.025 \
 U0LEXP =0.95 \
 UA =0.4007 \
 UAW =0.05 \
 UAWEXP =1 \
 UAL =0.00475 \
 UALEXP =1.118 \
 EUW =-0.02 \
 EUWEXP =1 \
 EUL =0.001 \
 EULEXP =1 \
 EU =1.9 \
 UDL =1E-15 \
 UDLEXP =1 \
 UD =1.042E-05 \
 UCS =2 \
 UCW =0 \
 UCWEXP =1 \
 UC =1E-07 \
 UCL =2.5E+04 \
 UCLEXP =1 \
 PCLM =0.15 \
 PCLML =0.01 \
 PCLMLEXP =0.4 \
 PCLMG =0 \
 PSCBE1 =5 \
 PSCBE2 =1.29E-12 \
 PDITS =0 \
 PDITSL =0 \
 PDITSD =0 \
 RSWMIN =0 \
 RSW =100 \
 RDWMIN =0 \
 RDW =100 \
 RDSW =20 \
 RDSWMIN =0 \
 PRWG =1 \
 PRWB =0 \
 WR =1 \
 RSH =0 \
 PDIBLCB =0 \
 PDIBLC =0.01 \
 PDIBLCL =1E-05 \
 PDIBLCLEXP =1E-06 \
 PVAG =0 \
 PTWG =0.2 \
 PTWGL =3E+04 \
 PTWGLEXP =5E-06 \
 FPROUT =0 \
 CF =0 \
 CFRCOEFF =1 \
 CGSO =2.5E-10 \
 CGDO =2.5E-10 \
 CGSL =1.2E-10 \
 CGDL =1.2E-10 \
 CKAPPAS =1.25 \
 CKAPPAD =1.25 \
 CGBO =0 \
 ADOS =0 \
 BDOS =1 \
 QM0 =0.001 \
 ETAQM =0.54 \
 NDEPCV =8E+23 \
 VFBCV =-0.95 \
 VSATCV =1E+05 \
 PCLMCV =0 \
 PSAT =0.46 \
 PSATL =6 \
 PSATLEXP =0.06 \
 TNFACTOR =0 \
 TETA0 =0 \
 UTE =-1.4 \
 UTEL =-0.001 \
 UA1 =-0.0011 \
 UA1L =0 \
 UC1 =0 \
 UD1 =0 \
 UD1L =0 \
 UCSTE =-0.005 \
 PRT =0 \
 AT =-0.05 \
 ATL =-0.1 \
 TDELTA =-0.0048 \
 PTWGT =-0.002 \
 PTWGTL =0.01 \
 KT1 =-0.115 \
 KT1EXP =1 \
 KT1L =1.286E-09 \
 KT2 =-0.003157 \
 K2LEXP =1.698 \
 K2WEXP =0.005 \
 TBGASUB =0 \
 IGCMOD =0 \
 IGBMOD =0 \
 AIGS=0.0136 \
 BIGS=0.00171 \
 CIGS=0.075 \
 AIGSL=0 \
 AIGD=0.0136 \
 BIGD=0.00171 \
 CIGD=0.075 \
 AIGDL=0 \
 AIGC=0.01285 \
 LAIGC=2.132E-06 \
 BIGC=0.0013 \
 CIGC=0.013 \
 AIGCL=-0.01227 \
 PIGCD=1 \
 PIGCDL=6.196 \
 AIGBINV=0.015 \
 BIGBINV=0.000949 \
 CIGBINV=0.006 \
 EIGBINV=1.1 \
 NIGBINV=3 \
 AIGBACC=0.01751 \
 BIGBACC=8.307 \
 CIGBACC=-898.7 \
 NIGBACC=1 \
 LPSAT=0 \
 WPSAT=0 \
 PPSAT=0 \
 PSATB=0 \
 PSATX=3 \
 WVSAT=0 \
 PVSAT=0 \
 WPTWG=0 \
 PPTWG=0 \
 TNOM=25 \
 WDVTP0=0 \
 WDVTP1=0 \
 LUTE=0.04574 \
 LUA1=8.365E-05 \
 LAT=0 \
 DVTP2=0 \
 DVTP3=0 \
 DVTP4=0 \
 DVTP5=0 \
 VSATL=1350 \
 VSATLEXP=0.00033 \
 SHMOD = 0 \
 RTH0 = 10m \
 MOBSCALE = 1
    

M_B (D G 0 0) bsim

simulator lang = spice

VD D  0 DC 1

simulator lang = spectre

VG (G  0) vsource dc=0.8 type=sine freq=1M sinedc=0.5 ampl=0.4

tranana tran start=0s stop=50ns step=00.0001ns maxstep=0.0001ns minstep=0.0001ns save=nooutput 






