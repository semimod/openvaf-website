Cir

.options reltol=1e-6 vabstol=1e-6 iabstol=1e-12 temp=26.85 save=nooutput

simulator lang = spectre


; Netlist

model bsim bsimsoi type=n version=4.4 \
 binunit = (1)             \
 mobmod  = (1)             \
 capmod  = (3)             \
 shmod   = (0)             \
 paramchk= (0)             \
 soimod  = (0)             \
 igcmod  = (1)             \
 igbmod  = (1)             \
 tsi     = (9e-008)        \
 tox     = (2e-009)        \
 toxref  = (2e-009)        \
 tbox    = (4e-007)        \
 toxqm   = (2e-009)        \
 tnom    = (27)            \
 rbody   = (0)             \
 rbsh    = (0)             \
 rsh     = (0)             \
 dtoxcv  = (0)             \
 xj      = (7e-008)        \
 rhalo   = (0)             \
 nch     = (1e+019)        \
 ngate   = (3e+020)        \
 wint    = (5.5544e-009)   \
 lint    = (2e-009)        \
 xpart   = (1)             \
 toxm    = (2e-009)        \
 k1      = (0.6)           \
 k2      = (1e-010)        \
 k3      = (0.231)         \
 k3b     = (0)             \
 kb1     = (1)             \
 w0      = (0)             \
 dvt0    = (2.2)           \
 dvt1    = (0.53)          \
 dvt2    = (0.127)         \
 dvt0w   = (0)             \
 dvt1w   = (0)             \
 dvt2w   = (0)             \
 eta0    = (1.7958)        \
 etab    = (-0.07)         \
 dsub    = (1.7577)        \
 voff    = (-0.10382)      \
 nfactor = (1)             \
 cdsc    = (0.00024)       \
 cdscb   = (0)             \
 cdscd   = (0)             \
 cit     = (0)             \
 u0      = (200)           \
 ua      = (2.25e-009)     \
 ub      = (5.9e-019)      \
 uc      = (2.9e-011)      \
 prwg    = (2.5)           \
 prwb    = (0.76)          \
 wr      = (1)             \
 rdsw    = (0.695)         \
 a0      = (0)             \
 ags     = (0)             \
 a1      = (0)             \
 a2      = (0.7)           \
 b0      = (0)             \
 b1      = (0)             \
 vsat    = (99820)         \
 keta    = (0)             \
 ketas   = (0)             \
 dwg     = (0)             \
 dwb     = (0)             \
 dwbc    = (0)             \
 pclm    = (1.3)           \
 pdiblc1 = (0.39)          \
 pdiblc2 = (0.05)          \
 pdiblcb = (0.89459)       \
 drout   = (2)             \
 pvag    = (0.116)         \
 delta   = (0.01)          \
 vevb    = (0.075)         \
 vecb    = (0.026)         \
 alpha0  = (5.0707e-009)   \
 beta0   = (0.0007605)     \
 beta1   = (0.0002767)     \
 beta2   = (0.094512)      \
 alphagb1= (0.35)          \
 alphagb2= (0.43)          \
 betagb1 = (0.03)          \
 betagb2 = (0.05)          \
 fbjtii  = (0)             \
 vdsatii0= (0.72051)       \
 tii     = (-0.5062)       \
 lii     = (2.835e-009)    \
 esatii  = (2213500)       \
 sii0    = (2.0387)        \
 sii1    = (0.04093)       \
 sii2    = (9.8e-011)      \
 siid    = (0.008025)      \
 aigc    = (1)             \
 bigc    = (0.05022)       \
 cigc    = (0.075)         \
 aigsd   = (0.43)          \
 bigsd   = (0.054)         \
 cigsd   = (0.075)         \
 nigc    = (1)             \
 poxedge = (1)             \
 pigcd   = (1)             \
 agidl   = (0)             \
 bgidl   = (0)             \
 ebg     = (1.2)           \
 vgb1    = (300)           \
 vgb2    = (17)            \
 voxh    = (1.5)           \
 deltavox= (0.004)         \
 ntox    = (1)             \
 ntun    = (1)             \
 ndiode  = (1)             \
 nrecf0  = (1.5)           \
 nrecr0  = (2)             \
 isbjt   = (1e-006)        \
 isdif   = (0.0001)        \
 isrec   = (0.01)          \
 istun   = (5e-005)        \
 vrec0   = (1)             \
 vtun0   = (0)             \
 nbjt    = (0.7888)        \
 lbjt0   = (1.4381e-006)   \
 vabjt   = (0.001)         \
 aely    = (1.0819e+010)   \
 ahli    = (0)             \
 lpe0    = (3e-009)        \
 cjswg   = (1e-010)        \
 mjswg   = (0.5)           \
 pbswg   = (0.7)           \
 tt      = (4e-010)        \
 ldif0   = (1)             \
 cgso    = (5e-011)        \
 cgdo    = (5e-011)        \
 dlc     = (0)             \
 dwc     = (0)             \
 dlcb    = (0)             \
 dlbg    = (0)             \
 fbody   = (1)             \
 clc     = (1e-008)        \
 cle     = (0)             \
 cf      = (0)             \
 csdmin  = (0)             \
 asd     = (0.3)           \
 csdesw  = (8.73e-011)     \
 delvt   = (-0.031456)     \
 acde    = (1)             \
 moin    = (25)            \
 ckappa  = (3.2309)        \
 cgdl    = (1.5533e-010)   \
 cgsl    = (1.5533e-010)   \
 ndif    = (-1)            \
 kt1     = (-0.11573)      \
 kt1l    = (-4e-010)       \
 kt2     = (-0.25)         \
 ute     = (-1.2189)       \
 ua1     = (5.005e-012)    \
 ub1     = (-8.835e-019)   \
 uc1     = (-6e-011)       \
 prt     = (51.149)        \
 rth0    = (0.02)          \
 cth0    = (1e-005)        \
 at      = (8479)          \
 tpbswg  = (5.86e-005)     \
 tcjswg  = (0.00092578)    \
 ntrecf  = (-0.55338)      \
 ntrecr  = (-0.15688)      \
 xbjt    = (1.0968)        \
 xdif    = (1.4551)        \
 xrec    = (2.6e-011)      \
 xtun    = (25.308)        \
 fnoimod = (0)             \
 tnoimod = (2)             \
 af      = (2.15)          \
 ef      = (1.119)         \
 kf      = (1.67e-026)     \
 w0flk   = (0.001)    

M_B (D G 0 0) bsim

simulator lang = spice

VG G  0 DC 0
VD D  0 DC 0

simulator lang = spectre

*dc_analysis dc start=0 stop=2 step=0.001 dev=VC useprevic=yes save=nooutput print=yes ; 

swp_vds sweep dev=VG start=0.5 stop=0.8 step=0.001 {
   dc_analysis dc start=0 stop=2 step=0.001 dev=VD useprevic=yes save=nooutput print=yes ; 
}






