HICUM/L2 Output Characteristics Xyce Simulation
.options nonlin reltol=1e-6 abstol=1e-12
.options device temp=26.85

* Netlist
.model hic npn level=234
.INCLUDE "model.lib"

Qt n_C n_B 0 0 n_TNODE hic

.PARAM V_B=0
.PARAM V_C=0

VV_B n_B 0 DC {V_B} 
VV_C n_C 0 DC {V_C}

.DC V_C 0 2 0.001 V_B 0.65 0.9 0.001 

.PRINT DC V(n_B) V(n_C)


.END
