HICUM/L2 Output Characteristics Xyce Simulation
.options nonlin reltol=1e-6 abstol=1e-12
.options device temp=26.85

* Netlist
.INCLUDE "bsim_built_in.lib"

Mt n_D n_G 0 0 BSI

.PARAM V_G=0
.PARAM V_D=0

VV_G n_G 0 DC {V_G} 
VV_D n_D 0 DC {V_D}

.DC V_D 0 2 0.001 V_G 0.5 0.8 0.01 



.END
