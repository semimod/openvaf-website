DMT Xyce simulation

* Netlist
YhicumL2_test Q_H n_C n_B n_E n_S n_TNODE _0
.MODEL _0 hicumL2_test abet = 2.4000000000e+01 acbar = 1.5000000000e+00 af = 2.0000000000e+00 afre = 2.0000000000e+00 ahc = 5.0000000000e-02 ahjei = 3.0000000000e+00 aick = 1.0000000000e-03 ajei = 1.6500000000e+00 ajep = 1.6000000000e+00 alb = 0.0000000000e+00 alces = -2.2860000000e-01 alfav = -2.4000000000e-03 alit = 3.3333300000e-01 alkav = 0.0000000000e+00 alqav = -6.2840000000e-04 alqf = 1.6666700000e-01 alrth = 0.0000000000e+00 alt0 = 4.0000000000e-03 alvs = 1.0000000000e-03 c10 = 9.0740000000e-30 cbcpar = 1.6451200000e-14 cbepar = 2.6090000000e-14 cfbe = -1 cjci0 = 3.5800000000e-15 cjcx0 = 6.2990000000e-15 cjei0 = 8.8690000000e-15 cjep0 = 2.1780000000e-15 cjs0 = 2.6000000000e-14 cscp0 = 0.0000000000e+00 csu = 0.0000000000e+00 cth = 0.0000000000e+00 delck = 2.0000000000e+00 dt = 0.0000000000e+00 dt0h = 8.0000000000e-14 dvgbe = 0.0000000000e+00 f1vg = -1.0237700000e-04 f2vg = 4.3215000000e-04 favl = 1.8960000000e+01 fbcpar = 3.0000000000e-01 fbepar = 1.0000000000e+00 fcrbi = 0.0000000000e+00 fdqr0 = 0.0000000000e+00 fgeo = 7.4090000000e-01 flcomp = 2.3000000000e+00 flcono = 0 flnqs = 0 flsh = 0 fqi = 1.0000000000e+00 fthc = 7.0000000000e-01 gtfe = 3.5480000000e+00 hf0 = 4.0000000000e+01 hfc = 2.0040000000e+01 hfe = 1.0010000000e+01 hjci = 2.0000000000e-01 hjei = 3.3820000000e+00 ibcis = 4.6030000000e-17 ibcxs = 0.0000000000e+00 ibeis = 1.3280000000e-19 ibeps = 1.2600000000e-19 ibets = 0.0000000000e+00 icbar = 1.0000000000e-02 ich = 0.0000000000e+00 ireis = 1.5000000000e-14 ireps = 1.8000000000e-14 iscs = 0.0000000000e+00 itss = 0.0000000000e+00 kavl = 0.0000000000e+00 kf = 0.0000000000e+00 kfre = 0.0000000000e+00 kt0 = 6.5880000000e-05 latb = 0.0000000000e+00 latl = 0.0000000000e+00 mbci = 1.1500000000e+00 mbcx = 1.0000000000e+00 mbei = 1.0270000000e+00 mbep = 1.0420000000e+00 mcf = 1.0000000000e+00 mrei = 2.0000000000e+00 mrep = 1.8000000000e+00 msc = 1.0000000000e+00 msf = 1.0000000000e+00 qavl = 5.0920000000e-14 qp0 = 1.0080000000e-13 rbi0 = 4.4440000000e+00 rbx = 2.5680000000e+00 rci0 = 9.5230000000e+00 rcx = 2.4830000000e+00 re = 1.5110000000e+00 rhjei = 2.0000000000e+00 rsu = 0.0000000000e+00 rth = 0.0000000000e+00 t0 = 2.0890000000e-13 tbhrec = 1.0000000000e-10 tbvl = 8.2500000000e-14 tef0 = 3.2710000000e-13 thcs = 5.0010000000e-12 tnom = 2.6850000000e+01 tr = 0.0000000000e+00 tsf = 0.0000000000e+00 tunode = 1 type = 1 vcbar = 4.0000000000e-02 vces = 1.0000000000e-02 vdci = 8.2010000000e-01 vdcx = 8.2010000000e-01 vdei = 7.1400000000e-01 vdep = 8.5010000000e-01 vds = 9.9970000000e-01 vdsp = 6.0000000000e-01 vgb = 9.1000000000e-01 vgc = 1.1700000000e+00 vge = 1.1700000000e+00 vgs = 1.1700000000e+00 vlim = 6.9990000000e-01 vpt = 2.0000000000e+00 vptci = 1.7900000000e+00 vptcx = 1.9770000000e+00 vpts = 1.0000000000e+02 vptsp = 1.0000000000e+02 zci = 2.8570000000e-01 zcx = 2.8630000000e-01 zei = 2.4890000000e-01 zep = 2.6320000000e-01 zetabet = 4.8920000000e+00 zetaci = 5.8000000000e-01 zetact = 5.0000000000e+00 zetacx = 0.0000000000e+00 zetahjei = -5.0000000000e-01 zetarbi = 3.0020000000e-01 zetarbx = 6.0110000000e-02 zetarcx = -2.7680000000e-02 zetare = -9.6050000000e-01 zetarth = 0.0000000000e+00 zetavgbe = 7.0000000000e-01 zs = 4.2950000000e-01 zsp = 5.0000000000e-01
RRbm n_B_FORCED n_B R=0.001  
RI_B n_BX n_B_FORCED R=0 
CCbm n_B_FORCED n_B C=1  
RI_C n_CX n_C_FORCED R=0 
RRcm n_C_FORCED n_C R=0.001  
CCcm n_C_FORCED n_C C=1  
RI_E n_EX n_E_FORCED R=0 
RRem n_E_FORCED n_E R=0.001  
CCem n_E_FORCED n_E C=1  
VV_B n_BX 0 DC {V_B} AC 1V 0.0 
VV_C n_CX 0 DC {V_C} AC 1V 0.0 
VV_E n_EX 0 DC {V_E} AC 1V 0.0 
RI_S n_SX n_S R=0 
RR_S n_SX n_EX R=5  
RR_t n_TNODE 0 R=1e9  
.PARAM V_B=0
.PARAM V_C=0
.PARAM V_S=0
.PARAM V_E=0
.PARAM ac_switch=0
.PARAM V_B_ac=1-ac_switch
.PARAM V_C_ac=ac_switch
.PARAM V_S_ac=0
.PARAM V_E_ac=0

* Table of operation points and temperatures: 
.DATA TAB_SIMS
+  V_E  V_B  ac_switch  V_C  TEMP
+  0.0  0.0        0.0  0.0 26.85
+  0.0  0.0        1.0  0.0 26.85
+  0.0  0.1        0.0  0.1 26.85
+  0.0  0.1        1.0  0.1 26.85
+  0.0  0.2        0.0  0.2 26.85
+  0.0  0.2        1.0  0.2 26.85
+  0.0  0.3        0.0  0.3 26.85
+  0.0  0.3        1.0  0.3 26.85
+  0.0  0.4        0.0  0.4 26.85
+  0.0  0.4        1.0  0.4 26.85
+  0.0  0.5        0.0  0.5 26.85
+  0.0  0.5        1.0  0.5 26.85
+  0.0  0.6        0.0  0.6 26.85
+  0.0  0.6        1.0  0.6 26.85
+  0.0  0.7        0.0  0.7 26.85
+  0.0  0.7        1.0  0.7 26.85
+  0.0  0.8        0.0  0.8 26.85
+  0.0  0.8        1.0  0.8 26.85
+  0.0  0.9        0.0  0.9 26.85
+  0.0  0.9        1.0  0.9 26.85
+  0.0  1.0        0.0  1.0 26.85
+  0.0  1.0        1.0  1.0 26.85
.ENDDATA

* step through ops simulation
.STEP DATA=TAB_SIMS
* DC OP simulation
.OP 
* DC OP output definition
.PRINT AC_IC FORMAT=CSV FILE=DC.csv TEMP V(*) I(*) ac_switch 
* AC simulation
.AC DATA=TAB_FREQUENCIES 
.DATA TAB_FREQUENCIES 
+ FREQ 
+ 1e+08 1e+09 
.ENDDATA 
* AC output definition
.PRINT AC FORMAT=CSV FILE=AC.csv V(*) I(*) 

.END
