Options ASCII_Rawfile=no DuplicateFunc="warning" DuplicateParam="warning" I_AbsTol=1e-12 A I_RelTol=1e-6 ResourceUsage=yes Temp=26.850000000000023 UseNutmegFormat=yes V_AbsTol=1e-6 V V_RelTol=1e-6 

simulator lang = spectre

model hic bht version=2.40 updatelevel=3.0 \ 
 c10 =  9.074e-030  \ 
 qp0 =  1.008e-013  \ 
 hfe =  10.01  \ 
 hfc =  20.04  \ 
 hjei =  3.382  \
 hjci =  0.2  \
 ibeis =  1.328e-019  \
 mbei =  1.027  \
 ireis =  1.5e-014  \
 mrei =  2  \
 ibeps =  1.26e-019  \
 mbep =  1.042  \
 ireps =  1.8e-014  \
 mrep =  1.8  \
 mcf =  1  \
 tbhrec =  1e-010  \
 ibcis =  4.603e-017  \
 mbci =  1.15  \
 ibcxs =  0  \
 mbcx =  1  \
 ibets =  0.02035  \
 abet =  24  \
 tunode =  1  \
 favl =  18.96  \
 qavl =  5.092e-014  \
 alfav =  -0.0024  \
 alqav =  -0.0006284  \
 rbi0 =  4.444  \
 rbx =  2.568  \
 fgeo =  0.7409  \
 fdqr0 =  0  \
 fcrbi =  0  \
 fqi =  1  \
 re =  1.511  \
 rcx =  2.483  \
 itss =  0  \
 msf =  1  \
 iscs =  0  \
 msc =  1  \
 tsf =  0  \
 rsu =  0  \
 csu =  0  \
 cjei0 =  8.869e-015  \
 vdei =  0.714  \
 zei =  0.2489  \
 ajei =  1.65  \
 cjep0 =  2.178e-015  \
 vdep =  0.8501  \
 zep =  0.2632  \
 ajep =  1.6  \
 cjci0 =  3.58e-015  \
 vdci =  0.8201  \
 zci =  0.2857  \
 vptci =  1.79  \
 cjcx0 =  6.299e-015  \
 vdcx =  0.8201  \
 zcx =  0.2863  \
 vptcx =  1.977  \
 fbcpar =  0.3  \
 fbepar =  1  \
 cjs0 =  2.6e-014  \
 vds =  0.9997  \
 zs =  0.4295  \
 vpts =  100  \
 t0 =  2.089e-013  \
 dt0h =  8e-014  \
 tbvl =  8.25e-014  \
 tef0 =  3.271e-013  \
 gtfe =  3.548  \
 thcs =  5.001e-012  \
 ahc =  0.05  \
 fthc =  0.7  \
 rci0 =  9.523  \
 vlim =  0.6999  \
 vces =  0.01  \
 vpt =  2  \
 tr =  0  \
 cbepar =  2.609e-014  \
 cbcpar =  1.64512e-014  \
 alqf =  0.166667  \
 alit =  0.333333  \
 flnqs =  0  \
 kf =  0  \
 af =  2  \
 cfbe =  -1  \
 latb =  0  \
 latl =  0  \
 vgb =  0.91  \
 alt0 =  0.004  \
 kt0 =  6.588e-005  \
 zetaci =  0.58  \
 alvs =  0.001  \
 alces =  -0.2286  \
 zetarbi =  0.3002  \
 zetarbx =  0.06011  \
 zetarcx =  -0.02768  \
 zetare =  -0.9605  \
 zetacx =  0  \
 vge =  1.17  \
 vgc =  1.17  \
 vgs =  1.17  \
 f1vg =  -0.000102377  \
 f2vg =  0.00043215  \
 zetact =  5  \
 zetabet =  4.892  \
 flsh =  1  \
 rth =  1113.4  \
 cth =  6.841e-012  \
 zetarth =  0  \
 alrth =  0.002  \
 flcomp =  2.3  \
 tnom =  26.85  \
 dt =  0  \
 acbar =  1.5  \
 flcono =  0  \
 icbar =  0.01  \
 vcbar =  0.04  \
 zetavgbe =  0.7  \
 hf0 =  40  \
 ahjei =  3  \
 rhjei =  2  \
 delck =  2  \
 zetahjei =  -0.5  

Q_H (C B  0  0) hic 


V_B (B 0) vsource dc=V_B type=dc 
V_C (C 0) vsource dc=V_C type=dc 

parameters V_B=0
parameters V_C=0

simulator lang = ads


ParamSweep:Sweep1 SimInstanceName[1]="DC1" StatusLevel=2 SweepVar="V_C" SweepPlan="Sweep1_stim" 
SweepPlan: Sweep1_stim Start=0 Stop=2 Step=0.01 

DC:DC1 StatusLevel=2 DevOpPtLevel=0 UseFiniteDiff=no PrintOpPoint=no Restart=0 \

ParamSweep:Sweep2 SimInstanceName[1]="Sweep1" StatusLevel=2 SweepVar="V_B" SweepPlan="Sweep2_stim" 
SweepPlan: Sweep2_stim Start=0.65 Stop=0.9 Step=0.001 
