Options ASCII_Rawfile=no DuplicateFunc="warning" DuplicateParam="warning" I_AbsTol=1e-12 A I_RelTol=1e-6 ResourceUsage=yes Temp=26.850000000000023 UseNutmegFormat=yes V_AbsTol=1e-6 V V_RelTol=1e-6 

#load "veriloga", "psp103.va"

; Netlist
PSP103VA:Q_H 0  0  0 0
R:Rb n_B 0 R=1e3

V_Source:V_B n_B 0 Vdc=V_B 

V_B=0

; simulation controllers
DC:DC SweepVar="V_B" SweepPlan="V_B_Plan" StatusLevel=0 DevOpPtLevel=4

; sweep plans
SweepPlan:V_B_Plan Start=0 Stop=0.01 Step=2



